`define ADD 6'h00
`define SUB 6'h01
`define MUL 6'h02
`define LDB 6'h10
`define LDW 6'h11
`define STB 6'h12
`define STW 6'h13
`define MOV 6'h14
`define BEQ 6'h30
`define JUMP 6'h31
`define TLBWRITE 6'h32
`define IRET 6'h33

`define ALU_X 31'hxxxxxxxx
