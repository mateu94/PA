`define ADD 7'h00
`define SUB 7'h01
`define MUL 7'h02
`define LDB 7'h10
`define LDW 7'h11
`define STB 7'h12
`define STW 7'h13
`define MOV 7'h14
`define BEQ 7'h30
`define JUMP 7'h31
`define TLBWRITE 7'h32
`define IRET 7'h33
`define X32 32'hXXXXXXXX